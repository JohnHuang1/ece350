module moduleName #(
    parameter N=2
) (
    input [N-1:0] a, b,
    input eq_prev, gt_prev,
    output eq, gt
);

    

endmodule