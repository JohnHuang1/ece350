// module moduleName #(
//     parameter N=32
// ) (
//     input[N-1:0] a, b,
//     output isEqual, isGreater
// );
//     // isEqual = a == b
//     // isGreater = a > b

    
    
// endmodule